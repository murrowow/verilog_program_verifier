module formula(a, b, out);
	input [1:0] a, b;
	output [1:0] cout;

	assign cout = a + b; 

endmodule
